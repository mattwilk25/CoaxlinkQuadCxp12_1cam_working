module udivision_LUT_8bit_int_to_64bit_frac #(
)(
    input logic [8-1:0] number_in,
    output logic [64-1:0] reciprocal

);

    logic [2**8-1:0] reciprocal_LUT [64-1:0];

    always_comb begin
        case (number_in)
        8'b00000000 : reciprocal = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        8'b00000001 : reciprocal = 64'b1000000000000000000000000000000000000000000000000000000000000000;
        8'b00000010 : reciprocal = 64'b0101010101010101010101010101010101010101010101010101010000000000;
        8'b00000011 : reciprocal = 64'b0100000000000000000000000000000000000000000000000000000000000000;
        8'b00000100 : reciprocal = 64'b0011001100110011001100110011001100110011001100110011010000000000;
        8'b00000101 : reciprocal = 64'b0010101010101010101010101010101010101010101010101010101000000000;
        8'b00000110 : reciprocal = 64'b0010010010010010010010010010010010010010010010010010010000000000;
        8'b00000111 : reciprocal = 64'b0010000000000000000000000000000000000000000000000000000000000000;
        8'b00001000 : reciprocal = 64'b0001110001110001110001110001110001110001110001110001110000000000;
        8'b00001001 : reciprocal = 64'b0001100110011001100110011001100110011001100110011001101000000000;
        8'b00001010 : reciprocal = 64'b0001011101000101110100010111010001011101000101110100011000000000;
        8'b00001011 : reciprocal = 64'b0001010101010101010101010101010101010101010101010101010100000000;
        8'b00001100 : reciprocal = 64'b0001001110110001001110110001001110110001001110110001010000000000;
        8'b00001101 : reciprocal = 64'b0001001001001001001001001001001001001001001001001001001000000000;
        8'b00001110 : reciprocal = 64'b0001000100010001000100010001000100010001000100010001000100000000;
        8'b00001111 : reciprocal = 64'b0001000000000000000000000000000000000000000000000000000000000000;
        8'b00010000 : reciprocal = 64'b0000111100001111000011110000111100001111000011110000111100000000;
        8'b00010001 : reciprocal = 64'b0000111000111000111000111000111000111000111000111000111000000000;
        8'b00010010 : reciprocal = 64'b0000110101111001010000110101111001010000110101111001010000000000;
        8'b00010011 : reciprocal = 64'b0000110011001100110011001100110011001100110011001100110100000000;
        8'b00010100 : reciprocal = 64'b0000110000110000110000110000110000110000110000110000110000000000;
        8'b00010101 : reciprocal = 64'b0000101110100010111010001011101000101110100010111010001100000000;
        8'b00010110 : reciprocal = 64'b0000101100100001011001000010110010000101100100001011001000000000;
        8'b00010111 : reciprocal = 64'b0000101010101010101010101010101010101010101010101010101010000000;
        8'b00011000 : reciprocal = 64'b0000101000111101011100001010001111010111000010100011110110000000;
        8'b00011001 : reciprocal = 64'b0000100111011000100111011000100111011000100111011000101000000000;
        8'b00011010 : reciprocal = 64'b0000100101111011010000100101111011010000100101111011010000000000;
        8'b00011011 : reciprocal = 64'b0000100100100100100100100100100100100100100100100100100100000000;
        8'b00011100 : reciprocal = 64'b0000100011010011110111001011000010001101001111011100101100000000;
        8'b00011101 : reciprocal = 64'b0000100010001000100010001000100010001000100010001000100010000000;
        8'b00011110 : reciprocal = 64'b0000100001000010000100001000010000100001000010000100001000000000;
        8'b00011111 : reciprocal = 64'b0000100000000000000000000000000000000000000000000000000000000000;
        8'b00100000 : reciprocal = 64'b0000011111000001111100000111110000011111000001111100001000000000;
        8'b00100001 : reciprocal = 64'b0000011110000111100001111000011110000111100001111000011110000000;
        8'b00100010 : reciprocal = 64'b0000011101010000011101010000011101010000011101010000011101000000;
        8'b00100011 : reciprocal = 64'b0000011100011100011100011100011100011100011100011100011100000000;
        8'b00100100 : reciprocal = 64'b0000011011101011001111100100010100110000011011101011010000000000;
        8'b00100101 : reciprocal = 64'b0000011010111100101000011010111100101000011010111100101000000000;
        8'b00100110 : reciprocal = 64'b0000011010010000011010010000011010010000011010010000011010000000;
        8'b00100111 : reciprocal = 64'b0000011001100110011001100110011001100110011001100110011010000000;
        8'b00101000 : reciprocal = 64'b0000011000111110011100000110001111100111000001100011111010000000;
        8'b00101001 : reciprocal = 64'b0000011000011000011000011000011000011000011000011000011000000000;
        8'b00101010 : reciprocal = 64'b0000010111110100000101111101000001011111010000010111110100000000;
        8'b00101011 : reciprocal = 64'b0000010111010001011101000101110100010111010001011101000110000000;
        8'b00101100 : reciprocal = 64'b0000010110110000010110110000010110110000010110110000010111000000;
        8'b00101101 : reciprocal = 64'b0000010110010000101100100001011001000010110010000101100100000000;
        8'b00101110 : reciprocal = 64'b0000010101110010011000100000101011100100110001000001010111000000;
        8'b00101111 : reciprocal = 64'b0000010101010101010101010101010101010101010101010101010101000000;
        8'b00110000 : reciprocal = 64'b0000010100111001011110000010100111001011110000010100111001000000;
        8'b00110001 : reciprocal = 64'b0000010100011110101110000101000111101011100001010001111011000000;
        8'b00110010 : reciprocal = 64'b0000010100000101000001010000010100000101000001010000010100000000;
        8'b00110011 : reciprocal = 64'b0000010011101100010011101100010011101100010011101100010100000000;
        8'b00110100 : reciprocal = 64'b0000010011010100100001110011111011001010110111100011000001000000;
        8'b00110101 : reciprocal = 64'b0000010010111101101000010010111101101000010010111101101000000000;
        8'b00110110 : reciprocal = 64'b0000010010100111100100000100101001111001000001001010011110000000;
        8'b00110111 : reciprocal = 64'b0000010010010010010010010010010010010010010010010010010010000000;
        8'b00111000 : reciprocal = 64'b0000010001111101110000010001111101110000010001111101110000000000;
        8'b00111001 : reciprocal = 64'b0000010001101001111011100101100001000110100111101110010110000000;
        8'b00111010 : reciprocal = 64'b0000010001010110110001111001011111011101010010011100001101000000;
        8'b00111011 : reciprocal = 64'b0000010001000100010001000100010001000100010001000100010001000000;
        8'b00111100 : reciprocal = 64'b0000010000110010010111000101001111101111001101101000111011000000;
        8'b00111101 : reciprocal = 64'b0000010000100001000010000100001000010000100001000010000100000000;
        8'b00111110 : reciprocal = 64'b0000010000010000010000010000010000010000010000010000010000000000;
        8'b00111111 : reciprocal = 64'b0000010000000000000000000000000000000000000000000000000000000000;
        8'b01000000 : reciprocal = 64'b0000001111110000001111110000001111110000001111110000010000000000;
        8'b01000001 : reciprocal = 64'b0000001111100000111110000011111000001111100000111110000100000000;
        8'b01000010 : reciprocal = 64'b0000001111010010001001100011010101111110000101101110110011100000;
        8'b01000011 : reciprocal = 64'b0000001111000011110000111100001111000011110000111100001111000000;
        8'b01000100 : reciprocal = 64'b0000001110110101110011000000111011010111001100000011101101100000;
        8'b01000101 : reciprocal = 64'b0000001110101000001110101000001110101000001110101000001110100000;
        8'b01000110 : reciprocal = 64'b0000001110011011000010101101000100100000011100110110000101100000;
        8'b01000111 : reciprocal = 64'b0000001110001110001110001110001110001110001110001110001110000000;
        8'b01001000 : reciprocal = 64'b0000001110000001110000001110000001110000001110000001110000000000;
        8'b01001001 : reciprocal = 64'b0000001101110101100111110010001010011000001101110101101000000000;
        8'b01001010 : reciprocal = 64'b0000001101101001110100000011011010011101000000110110100111100000;
        8'b01001011 : reciprocal = 64'b0000001101011110010100001101011110010100001101011110010100000000;
        8'b01001100 : reciprocal = 64'b0000001101010011000111011110110000001101010011000111011111000000;
        8'b01001101 : reciprocal = 64'b0000001101001000001101001000001101001000001101001000001101000000;
        8'b01001110 : reciprocal = 64'b0000001100111101100100011101001010100010000001100111101100100000;
        8'b01001111 : reciprocal = 64'b0000001100110011001100110011001100110011001100110011001101000000;
        8'b01010000 : reciprocal = 64'b0000001100101001000101100001111110011010110111010011110000000000;
        8'b01010001 : reciprocal = 64'b0000001100011111001110000011000111110011100000110001111101000000;
        8'b01010010 : reciprocal = 64'b0000001100010101100101110010000111101101011111100111010101000000;
        8'b01010011 : reciprocal = 64'b0000001100001100001100001100001100001100001100001100001100000000;
        8'b01010100 : reciprocal = 64'b0000001100000011000000110000001100000011000000110000001100000000;
        8'b01010101 : reciprocal = 64'b0000001011111010000010111110100000101111101000001011111010000000;
        8'b01010110 : reciprocal = 64'b0000001011110001010010011001000000101111000101001001100100000000;
        8'b01010111 : reciprocal = 64'b0000001011101000101110100010111010001011101000101110100011000000;
        8'b01011000 : reciprocal = 64'b0000001011100000010111000000101110000001011100000010111000000000;
        8'b01011001 : reciprocal = 64'b0000001011011000001011011000001011011000001011011000001011100000;
        8'b01011010 : reciprocal = 64'b0000001011010000001011010000001011010000001011010000001011100000;
        8'b01011011 : reciprocal = 64'b0000001011001000010110010000101100100001011001000010110010000000;
        8'b01011100 : reciprocal = 64'b0000001011000000101100000010110000001011000000101100000011000000;
        8'b01011101 : reciprocal = 64'b0000001010111001001100010000010101110010011000100000101011100000;
        8'b01011110 : reciprocal = 64'b0000001010110001110110100100011000010000001010110001110110100000;
        8'b01011111 : reciprocal = 64'b0000001010101010101010101010101010101010101010101010101010100000;
        8'b01100000 : reciprocal = 64'b0000001010100011101000001111110101011100010111110000001010100000;
        8'b01100001 : reciprocal = 64'b0000001010011100101111000001010011100101111000001010011100100000;
        8'b01100010 : reciprocal = 64'b0000001010010101111110101101010000001010010101111110101101100000;
        8'b01100011 : reciprocal = 64'b0000001010001111010111000010100011110101110000101000111101100000;
        8'b01100100 : reciprocal = 64'b0000001010001000110111110000110010101100010110110011111101100000;
        8'b01100101 : reciprocal = 64'b0000001010000010100000101000001010000010100000101000001010000000;
        8'b01100110 : reciprocal = 64'b0000001001111100010001011001011110011100100101010010000001000000;
        8'b01100111 : reciprocal = 64'b0000001001110110001001110110001001110110001001110110001010000000;
        8'b01101000 : reciprocal = 64'b0000001001110000001001110000001001110000001001110000001010000000;
        8'b01101001 : reciprocal = 64'b0000001001101010010000111001111101100101011011110001100000100000;
        8'b01101010 : reciprocal = 64'b0000001001100100011111000110100101000101011000100001011111100000;
        8'b01101011 : reciprocal = 64'b0000001001011110110100001001011110110100001001011110110100000000;
        8'b01101100 : reciprocal = 64'b0000001001011001001111110110100110110000001001011001010000000000;
        8'b01101101 : reciprocal = 64'b0000001001010011110010000010010100111100100000100101001111000000;
        8'b01101110 : reciprocal = 64'b0000001001001110011010100001011100010000001001001110011010100000;
        8'b01101111 : reciprocal = 64'b0000001001001001001001001001001001001001001001001001001001000000;
        8'b01110000 : reciprocal = 64'b0000001001000011111101101111000000100100001111110110111100000000;
        8'b01110001 : reciprocal = 64'b0000001000111110111000001000111110111000001000111110111000000000;
        8'b01110010 : reciprocal = 64'b0000001000111001111000001101010110110100010100000010001110100000;
        8'b01110011 : reciprocal = 64'b0000001000110100111101110010110000100011010011110111001011000000;
        8'b01110100 : reciprocal = 64'b0000001000110000001000110000001000110000001000110000001001000000;
        8'b01110101 : reciprocal = 64'b0000001000101011011000111100101111101110101001001110000110100000;
        8'b01110110 : reciprocal = 64'b0000001000100110101110010000001000100110101110010000001000100000;
        8'b01110111 : reciprocal = 64'b0000001000100010001000100010001000100010001000100010001000100000;
        8'b01111000 : reciprocal = 64'b0000001000011101100111101010110101111100110100111001001000000000;
        8'b01111001 : reciprocal = 64'b0000001000011001001011100010100111110111100110110100011101100000;
        8'b01111010 : reciprocal = 64'b0000001000010100110100000010000101001101000000100001010011100000;
        8'b01111011 : reciprocal = 64'b0000001000010000100001000010000100001000010000100001000010000000;
        8'b01111100 : reciprocal = 64'b0000001000001100010010011011101001011110001101010011111110000000;
        8'b01111101 : reciprocal = 64'b0000001000001000001000001000001000001000001000001000001000000000;
        8'b01111110 : reciprocal = 64'b0000001000000100000010000001000000100000010000001000000100000000;
        8'b01111111 : reciprocal = 64'b0000001000000000000000000000000000000000000000000000000000000000;
        8'b10000000 : reciprocal = 64'b0000000111111100000001111111000000011111110000000111111100000000;
        8'b10000001 : reciprocal = 64'b0000000111111000000111111000000111111000000111111000001000000000;
        8'b10000010 : reciprocal = 64'b0000000111110100010001100101100111100100101001000010011100010000;
        8'b10000011 : reciprocal = 64'b0000000111110000011111000001111100000111110000011111000010000000;
        8'b10000100 : reciprocal = 64'b0000000111101100110000000111101100110000000111101100110000000000;
        8'b10000101 : reciprocal = 64'b0000000111101001000100110001101010111111000010110111011001110000;
        8'b10000110 : reciprocal = 64'b0000000111100101011100111010110010010000000111100101011101000000;
        8'b10000111 : reciprocal = 64'b0000000111100001111000011110000111100001111000011110000111100000;
        8'b10001000 : reciprocal = 64'b0000000111011110010111010110111000111111100010000110100010100000;
        8'b10001001 : reciprocal = 64'b0000000111011010111001100000011101101011100110000001110110110000;
        8'b10001010 : reciprocal = 64'b0000000111010111011110110110010101001011100000101100001101000000;
        8'b10001011 : reciprocal = 64'b0000000111010100000111010100000111010100000111010100000111010000;
        8'b10001100 : reciprocal = 64'b0000000111010000110010110101100011110110111011000000011101000000;
        8'b10001101 : reciprocal = 64'b0000000111001101100001010110100010010000001110011011000010110000;
        8'b10001110 : reciprocal = 64'b0000000111001010010010110011000001010101111011100001100100010000;
        8'b10001111 : reciprocal = 64'b0000000111000111000111000111000111000111000111000111000111000000;
        8'b10010000 : reciprocal = 64'b0000000111000011111110001111000000011100001111111000111100000000;
        8'b10010001 : reciprocal = 64'b0000000111000000111000000111000000111000000111000000111000000000;
        8'b10010010 : reciprocal = 64'b0000000110111101110100101011100010011001010000000110111101110000;
        8'b10010011 : reciprocal = 64'b0000000110111010110011111001000101001100000110111010110100000000;
        8'b10010100 : reciprocal = 64'b0000000110110111110101101100001111011101101000110011100010110000;
        8'b10010101 : reciprocal = 64'b0000000110110100111010000001101101001110100000011011010011110000;
        8'b10010110 : reciprocal = 64'b0000000110110010000000110110010000000110110010000000110110010000;
        8'b10010111 : reciprocal = 64'b0000000110101111001010000110101111001010000110101111001010000000;
        8'b10011000 : reciprocal = 64'b0000000110101100010101110000000110101100010101110000000110110000;
        8'b10011001 : reciprocal = 64'b0000000110101001100011101111011000000110101001100011101111100000;
        8'b10011010 : reciprocal = 64'b0000000110100110110100000001101001101101000000011010011011010000;
        8'b10011011 : reciprocal = 64'b0000000110100100000110100100000110100100000110100100000110100000;
        8'b10011100 : reciprocal = 64'b0000000110100001011011010011111110010111101001001011000000100000;
        8'b10011101 : reciprocal = 64'b0000000110011110110010001110100101010001000000110011110110010000;
        8'b10011110 : reciprocal = 64'b0000000110011100001011010001010011101110010010100001000000100000;
        8'b10011111 : reciprocal = 64'b0000000110011001100110011001100110011001100110011001100110100000;
        8'b10100000 : reciprocal = 64'b0000000110010111000011100100111110000000110010111000011100100000;
        8'b10100001 : reciprocal = 64'b0000000110010100100010110000111111001101011011101001111000000000;
        8'b10100010 : reciprocal = 64'b0000000110010010000011111011010010011101000011100010001010010000;
        8'b10100011 : reciprocal = 64'b0000000110001111100111000001100011111001110000011000111110100000;
        8'b10100100 : reciprocal = 64'b0000000110001101001100000001100011010011000000011000110100110000;
        8'b10100101 : reciprocal = 64'b0000000110001010110010111001000011110110101111110011101010100000;
        8'b10100110 : reciprocal = 64'b0000000110001000011011100101111100001010101110110000010010100000;
        8'b10100111 : reciprocal = 64'b0000000110000110000110000110000110000110000110000110000110000000;
        8'b10101000 : reciprocal = 64'b0000000110000011110010010111011110101011001010111110110111010000;
        8'b10101001 : reciprocal = 64'b0000000110000001100000011000000110000001100000011000000110000000;
        8'b10101010 : reciprocal = 64'b0000000101111111010000000101111111010000000101111111010000000000;
        8'b10101011 : reciprocal = 64'b0000000101111101000001011111010000010111110100000101111101000000;
        8'b10101100 : reciprocal = 64'b0000000101111010110100100010000010001110000011101100110000110000;
        8'b10101101 : reciprocal = 64'b0000000101111000101001001100100000010111100010100100110010000000;
        8'b10101110 : reciprocal = 64'b0000000101110110011111011100111001000011010010101001101100010000;
        8'b10101111 : reciprocal = 64'b0000000101110100010111010001011101000101110100010111010001100000;
        8'b10110000 : reciprocal = 64'b0000000101110010010000101000011111110100011011011110101111000000;
        8'b10110001 : reciprocal = 64'b0000000101110000001011100000010111000000101110000001011100000000;
        8'b10110010 : reciprocal = 64'b0000000101101110000111110111011010110100001100110111110001110000;
        8'b10110011 : reciprocal = 64'b0000000101101100000101101100000101101100000101101100000101110000;
        8'b10110100 : reciprocal = 64'b0000000101101010000100111100110100010101001101110010100100000000;
        8'b10110101 : reciprocal = 64'b0000000101101000000101101000000101101000000101101000000101110000;
        8'b10110110 : reciprocal = 64'b0000000101100110000111101100011010100101000100100010111110010000;
        8'b10110111 : reciprocal = 64'b0000000101100100001011001000010110010000101100100001011001000000;
        8'b10111000 : reciprocal = 64'b0000000101100010001111111010011101110000000101100010010000000000;
        8'b10111001 : reciprocal = 64'b0000000101100000010110000001011000000101100000010110000001100000;
        8'b10111010 : reciprocal = 64'b0000000101011110011101011011101110001101000000010101111001110000;
        8'b10111011 : reciprocal = 64'b0000000101011100100110001000001010111001001100010000010101110000;
        8'b10111100 : reciprocal = 64'b0000000101011010110000000101011010110000000101011010110000000000;
        8'b10111101 : reciprocal = 64'b0000000101011000111011010010001100001000000101011000111011010000;
        8'b10111110 : reciprocal = 64'b0000000101010111000111101101001111000101000001101011001110100000;
        8'b10111111 : reciprocal = 64'b0000000101010101010101010101010101010101010101010101010101010000;
        8'b11000000 : reciprocal = 64'b0000000101010011100100001001010010001111010000001111111010110000;
        8'b11000001 : reciprocal = 64'b0000000101010001110100000111111010101110001011111000000101010000;
        8'b11000010 : reciprocal = 64'b0000000101010000000101010000000101010000000101010000000101010000;
        8'b11000011 : reciprocal = 64'b0000000101001110010111100000101001110010111100000101001110010000;
        8'b11000100 : reciprocal = 64'b0000000101001100101010111000100001110010010110101111011011100000;
        8'b11000101 : reciprocal = 64'b0000000101001010111111010110101000000101001010111111010110110000;
        8'b11000110 : reciprocal = 64'b0000000101001001010100111001111000111011001011010000011001110000;
        8'b11000111 : reciprocal = 64'b0000000101000111101011100001010001111010111000010100011110110000;
        8'b11001000 : reciprocal = 64'b0000000101000110000011001011110001111111010111001111100110100000;
        8'b11001001 : reciprocal = 64'b0000000101000100011011111000011001010110001011011001111110110000;
        8'b11001010 : reciprocal = 64'b0000000101000010110101100110001001011101010100011111100001110000;
        8'b11001011 : reciprocal = 64'b0000000101000001010000010100000101000001010000010100000101000000;
        8'b11001100 : reciprocal = 64'b0000000100111111101100000001001111111011000000010011111110110000;
        8'b11001101 : reciprocal = 64'b0000000100111110001000101100101111001110010010101001000000100000;
        8'b11001110 : reciprocal = 64'b0000000100111100100110010101101001000111101110101011111001110000;
        8'b11001111 : reciprocal = 64'b0000000100111011000100111011000100111011000100111011000101000000;
        8'b11010000 : reciprocal = 64'b0000000100111001100100011100001011000001100001111111011000110000;
        8'b11010001 : reciprocal = 64'b0000000100111000000100111000000100111000000100111000000101000000;
        8'b11010010 : reciprocal = 64'b0000000100110110100110001101111100111101111000000111010010000000;
        8'b11010011 : reciprocal = 64'b0000000100110101001000011100111110110010101101111000110000010000;
        8'b11010100 : reciprocal = 64'b0000000100110011101011100100010110110101011110111100101100100000;
        8'b11010101 : reciprocal = 64'b0000000100110010001111100011010010100010101100010000101111110000;
        8'b11010110 : reciprocal = 64'b0000000100110000110100011001000000010011000011010001100100000000;
        8'b11010111 : reciprocal = 64'b0000000100101111011010000100101111011010000100101111011010000000;
        8'b11011000 : reciprocal = 64'b0000000100101110000000100101110000000100101110000000100101110000;
        8'b11011001 : reciprocal = 64'b0000000100101100100111111011010011011000000100101100101000000000;
        8'b11011010 : reciprocal = 64'b0000000100101011010000000100101011010000000100101011010000000000;
        8'b11011011 : reciprocal = 64'b0000000100101001111001000001001010011110010000010010100111100000;
        8'b11011100 : reciprocal = 64'b0000000100101000100010110000000100101000100010110000000100110000;
        8'b11011101 : reciprocal = 64'b0000000100100111001101010000101110001000000100100111001101010000;
        8'b11011110 : reciprocal = 64'b0000000100100101111000100010011100001000000010010010111100010000;
        8'b11011111 : reciprocal = 64'b0000000100100100100100100100100100100100100100100100100100100000;
        8'b11100000 : reciprocal = 64'b0000000100100011010001010110011110001001101010111100110111110000;
        8'b11100001 : reciprocal = 64'b0000000100100001111110110111100000010010000111111011011110000000;
        8'b11100010 : reciprocal = 64'b0000000100100000101101000111000011000110011111000000110110010000;
        8'b11100011 : reciprocal = 64'b0000000100011111011100000100011111011100000100011111011100000000;
        8'b11100100 : reciprocal = 64'b0000000100011110001011101111001110110011111110111000011101000000;
        8'b11100101 : reciprocal = 64'b0000000100011100111100000110101011011010001010000001000111010000;
        8'b11100110 : reciprocal = 64'b0000000100011011101101001010010000000100011011101101001010010000;
        8'b11100111 : reciprocal = 64'b0000000100011010011110111001011000010001101001111011100101100000;
        8'b11101000 : reciprocal = 64'b0000000100011001010001010011100000001000110010100010100111000000;
        8'b11101001 : reciprocal = 64'b0000000100011000000100011000000100011000000100011000000100100000;
        8'b11101010 : reciprocal = 64'b0000000100010110111000000110100010010100001001110011011110010000;
        8'b11101011 : reciprocal = 64'b0000000100010101101100011110010111110111010100100111000011010000;
        8'b11101100 : reciprocal = 64'b0000000100010100100001011111000011100000101011001101001110110000;
        8'b11101101 : reciprocal = 64'b0000000100010011010111001000000100010011010111001000000100010000;
        8'b11101110 : reciprocal = 64'b0000000100010010001101011000111001110101110100110000001100110000;
        8'b11101111 : reciprocal = 64'b0000000100010001000100010001000100010001000100010001000100010000;
        8'b11110000 : reciprocal = 64'b0000000100001111111011110000000100001111111011110000000100010000;
        8'b11110001 : reciprocal = 64'b0000000100001110110011110101011010111110011010011100100100000000;
        8'b11110010 : reciprocal = 64'b0000000100001101101100100000101010001000111101000110100101100000;
        8'b11110011 : reciprocal = 64'b0000000100001100100101110001010011111011110011011010001110110000;
        8'b11110100 : reciprocal = 64'b0000000100001011011111100110111011000010010110011101110010000000;
        8'b11110101 : reciprocal = 64'b0000000100001010011010000001000010100110100000010000101001110000;
        8'b11110110 : reciprocal = 64'b0000000100001001010100111111001110010000000100001001010101000000;
        8'b11110111 : reciprocal = 64'b0000000100001000010000100001000010000100001000010000100001000000;
        8'b11111000 : reciprocal = 64'b0000000100000111001100100110000010100100011111110111110001100000;
        8'b11111001 : reciprocal = 64'b0000000100000110001001001101110100101111000110101001111111000000;
        8'b11111010 : reciprocal = 64'b0000000100000101000110010111111101111101011100110100000001000000;
        8'b11111011 : reciprocal = 64'b0000000100000100000100000100000100000100000100000100000100000000;
        8'b11111100 : reciprocal = 64'b0000000100000011000010010001101101010001111101011110000110100000;
        8'b11111101 : reciprocal = 64'b0000000100000010000001000000100000010000001000000100000010000000;
        8'b11111110 : reciprocal = 64'b0000000100000001000000010000000100000001000000010000000100000000;
        8'b11111111 : reciprocal = 64'b0000000100000000000000000000000000000000000000000000000000000000;


        endcase
    end
    



    //////////////////////// For testbenching ////////////////////////
    // synthesis translate_off

    // synthesis translate_on

endmodule
