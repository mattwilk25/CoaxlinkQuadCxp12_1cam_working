module udivision_LUT_8bit_int_to_16bit_frac #(
)(
    input logic [8-1:0] number_in,
    output logic [16-1:0] reciprocal

);

    logic [2**8-1:0] reciprocal_LUT [16-1:0];

    always_comb begin
        case (number_in)
        8'b00000000 : reciprocal = 16'b1111111111111111;
        8'b00000001 : reciprocal = 16'b1000000000000000;
        8'b00000010 : reciprocal = 16'b0101010101010101;
        8'b00000011 : reciprocal = 16'b0100000000000000;
        8'b00000100 : reciprocal = 16'b0011001100110011;
        8'b00000101 : reciprocal = 16'b0010101010101010;
        8'b00000110 : reciprocal = 16'b0010010010010010;
        8'b00000111 : reciprocal = 16'b0010000000000000;
        8'b00001000 : reciprocal = 16'b0001110001110001;
        8'b00001001 : reciprocal = 16'b0001100110011001;
        8'b00001010 : reciprocal = 16'b0001011101000101;
        8'b00001011 : reciprocal = 16'b0001010101010101;
        8'b00001100 : reciprocal = 16'b0001001110110001;
        8'b00001101 : reciprocal = 16'b0001001001001001;
        8'b00001110 : reciprocal = 16'b0001000100010001;
        8'b00001111 : reciprocal = 16'b0001000000000000;
        8'b00010000 : reciprocal = 16'b0000111100001111;
        8'b00010001 : reciprocal = 16'b0000111000111000;
        8'b00010010 : reciprocal = 16'b0000110101111001;
        8'b00010011 : reciprocal = 16'b0000110011001100;
        8'b00010100 : reciprocal = 16'b0000110000110000;
        8'b00010101 : reciprocal = 16'b0000101110100010;
        8'b00010110 : reciprocal = 16'b0000101100100001;
        8'b00010111 : reciprocal = 16'b0000101010101010;
        8'b00011000 : reciprocal = 16'b0000101000111101;
        8'b00011001 : reciprocal = 16'b0000100111011000;
        8'b00011010 : reciprocal = 16'b0000100101111011;
        8'b00011011 : reciprocal = 16'b0000100100100100;
        8'b00011100 : reciprocal = 16'b0000100011010011;
        8'b00011101 : reciprocal = 16'b0000100010001000;
        8'b00011110 : reciprocal = 16'b0000100001000010;
        8'b00011111 : reciprocal = 16'b0000100000000000;
        8'b00100000 : reciprocal = 16'b0000011111000001;
        8'b00100001 : reciprocal = 16'b0000011110000111;
        8'b00100010 : reciprocal = 16'b0000011101010000;
        8'b00100011 : reciprocal = 16'b0000011100011100;
        8'b00100100 : reciprocal = 16'b0000011011101011;
        8'b00100101 : reciprocal = 16'b0000011010111100;
        8'b00100110 : reciprocal = 16'b0000011010010000;
        8'b00100111 : reciprocal = 16'b0000011001100110;
        8'b00101000 : reciprocal = 16'b0000011000111110;
        8'b00101001 : reciprocal = 16'b0000011000011000;
        8'b00101010 : reciprocal = 16'b0000010111110100;
        8'b00101011 : reciprocal = 16'b0000010111010001;
        8'b00101100 : reciprocal = 16'b0000010110110000;
        8'b00101101 : reciprocal = 16'b0000010110010000;
        8'b00101110 : reciprocal = 16'b0000010101110010;
        8'b00101111 : reciprocal = 16'b0000010101010101;
        8'b00110000 : reciprocal = 16'b0000010100111001;
        8'b00110001 : reciprocal = 16'b0000010100011110;
        8'b00110010 : reciprocal = 16'b0000010100000101;
        8'b00110011 : reciprocal = 16'b0000010011101100;
        8'b00110100 : reciprocal = 16'b0000010011010100;
        8'b00110101 : reciprocal = 16'b0000010010111101;
        8'b00110110 : reciprocal = 16'b0000010010100111;
        8'b00110111 : reciprocal = 16'b0000010010010010;
        8'b00111000 : reciprocal = 16'b0000010001111101;
        8'b00111001 : reciprocal = 16'b0000010001101001;
        8'b00111010 : reciprocal = 16'b0000010001010110;
        8'b00111011 : reciprocal = 16'b0000010001000100;
        8'b00111100 : reciprocal = 16'b0000010000110010;
        8'b00111101 : reciprocal = 16'b0000010000100001;
        8'b00111110 : reciprocal = 16'b0000010000010000;
        8'b00111111 : reciprocal = 16'b0000010000000000;
        8'b01000000 : reciprocal = 16'b0000001111110000;
        8'b01000001 : reciprocal = 16'b0000001111100000;
        8'b01000010 : reciprocal = 16'b0000001111010010;
        8'b01000011 : reciprocal = 16'b0000001111000011;
        8'b01000100 : reciprocal = 16'b0000001110110101;
        8'b01000101 : reciprocal = 16'b0000001110101000;
        8'b01000110 : reciprocal = 16'b0000001110011011;
        8'b01000111 : reciprocal = 16'b0000001110001110;
        8'b01001000 : reciprocal = 16'b0000001110000001;
        8'b01001001 : reciprocal = 16'b0000001101110101;
        8'b01001010 : reciprocal = 16'b0000001101101001;
        8'b01001011 : reciprocal = 16'b0000001101011110;
        8'b01001100 : reciprocal = 16'b0000001101010011;
        8'b01001101 : reciprocal = 16'b0000001101001000;
        8'b01001110 : reciprocal = 16'b0000001100111101;
        8'b01001111 : reciprocal = 16'b0000001100110011;
        8'b01010000 : reciprocal = 16'b0000001100101001;
        8'b01010001 : reciprocal = 16'b0000001100011111;
        8'b01010010 : reciprocal = 16'b0000001100010101;
        8'b01010011 : reciprocal = 16'b0000001100001100;
        8'b01010100 : reciprocal = 16'b0000001100000011;
        8'b01010101 : reciprocal = 16'b0000001011111010;
        8'b01010110 : reciprocal = 16'b0000001011110001;
        8'b01010111 : reciprocal = 16'b0000001011101000;
        8'b01011000 : reciprocal = 16'b0000001011100000;
        8'b01011001 : reciprocal = 16'b0000001011011000;
        8'b01011010 : reciprocal = 16'b0000001011010000;
        8'b01011011 : reciprocal = 16'b0000001011001000;
        8'b01011100 : reciprocal = 16'b0000001011000000;
        8'b01011101 : reciprocal = 16'b0000001010111001;
        8'b01011110 : reciprocal = 16'b0000001010110001;
        8'b01011111 : reciprocal = 16'b0000001010101010;
        8'b01100000 : reciprocal = 16'b0000001010100011;
        8'b01100001 : reciprocal = 16'b0000001010011100;
        8'b01100010 : reciprocal = 16'b0000001010010101;
        8'b01100011 : reciprocal = 16'b0000001010001111;
        8'b01100100 : reciprocal = 16'b0000001010001000;
        8'b01100101 : reciprocal = 16'b0000001010000010;
        8'b01100110 : reciprocal = 16'b0000001001111100;
        8'b01100111 : reciprocal = 16'b0000001001110110;
        8'b01101000 : reciprocal = 16'b0000001001110000;
        8'b01101001 : reciprocal = 16'b0000001001101010;
        8'b01101010 : reciprocal = 16'b0000001001100100;
        8'b01101011 : reciprocal = 16'b0000001001011110;
        8'b01101100 : reciprocal = 16'b0000001001011001;
        8'b01101101 : reciprocal = 16'b0000001001010011;
        8'b01101110 : reciprocal = 16'b0000001001001110;
        8'b01101111 : reciprocal = 16'b0000001001001001;
        8'b01110000 : reciprocal = 16'b0000001001000011;
        8'b01110001 : reciprocal = 16'b0000001000111110;
        8'b01110010 : reciprocal = 16'b0000001000111001;
        8'b01110011 : reciprocal = 16'b0000001000110100;
        8'b01110100 : reciprocal = 16'b0000001000110000;
        8'b01110101 : reciprocal = 16'b0000001000101011;
        8'b01110110 : reciprocal = 16'b0000001000100110;
        8'b01110111 : reciprocal = 16'b0000001000100010;
        8'b01111000 : reciprocal = 16'b0000001000011101;
        8'b01111001 : reciprocal = 16'b0000001000011001;
        8'b01111010 : reciprocal = 16'b0000001000010100;
        8'b01111011 : reciprocal = 16'b0000001000010000;
        8'b01111100 : reciprocal = 16'b0000001000001100;
        8'b01111101 : reciprocal = 16'b0000001000001000;
        8'b01111110 : reciprocal = 16'b0000001000000100;
        8'b01111111 : reciprocal = 16'b0000001000000000;
        8'b10000000 : reciprocal = 16'b0000000111111100;
        8'b10000001 : reciprocal = 16'b0000000111111000;
        8'b10000010 : reciprocal = 16'b0000000111110100;
        8'b10000011 : reciprocal = 16'b0000000111110000;
        8'b10000100 : reciprocal = 16'b0000000111101100;
        8'b10000101 : reciprocal = 16'b0000000111101001;
        8'b10000110 : reciprocal = 16'b0000000111100101;
        8'b10000111 : reciprocal = 16'b0000000111100001;
        8'b10001000 : reciprocal = 16'b0000000111011110;
        8'b10001001 : reciprocal = 16'b0000000111011010;
        8'b10001010 : reciprocal = 16'b0000000111010111;
        8'b10001011 : reciprocal = 16'b0000000111010100;
        8'b10001100 : reciprocal = 16'b0000000111010000;
        8'b10001101 : reciprocal = 16'b0000000111001101;
        8'b10001110 : reciprocal = 16'b0000000111001010;
        8'b10001111 : reciprocal = 16'b0000000111000111;
        8'b10010000 : reciprocal = 16'b0000000111000011;
        8'b10010001 : reciprocal = 16'b0000000111000000;
        8'b10010010 : reciprocal = 16'b0000000110111101;
        8'b10010011 : reciprocal = 16'b0000000110111010;
        8'b10010100 : reciprocal = 16'b0000000110110111;
        8'b10010101 : reciprocal = 16'b0000000110110100;
        8'b10010110 : reciprocal = 16'b0000000110110010;
        8'b10010111 : reciprocal = 16'b0000000110101111;
        8'b10011000 : reciprocal = 16'b0000000110101100;
        8'b10011001 : reciprocal = 16'b0000000110101001;
        8'b10011010 : reciprocal = 16'b0000000110100110;
        8'b10011011 : reciprocal = 16'b0000000110100100;
        8'b10011100 : reciprocal = 16'b0000000110100001;
        8'b10011101 : reciprocal = 16'b0000000110011110;
        8'b10011110 : reciprocal = 16'b0000000110011100;
        8'b10011111 : reciprocal = 16'b0000000110011001;
        8'b10100000 : reciprocal = 16'b0000000110010111;
        8'b10100001 : reciprocal = 16'b0000000110010100;
        8'b10100010 : reciprocal = 16'b0000000110010010;
        8'b10100011 : reciprocal = 16'b0000000110001111;
        8'b10100100 : reciprocal = 16'b0000000110001101;
        8'b10100101 : reciprocal = 16'b0000000110001010;
        8'b10100110 : reciprocal = 16'b0000000110001000;
        8'b10100111 : reciprocal = 16'b0000000110000110;
        8'b10101000 : reciprocal = 16'b0000000110000011;
        8'b10101001 : reciprocal = 16'b0000000110000001;
        8'b10101010 : reciprocal = 16'b0000000101111111;
        8'b10101011 : reciprocal = 16'b0000000101111101;
        8'b10101100 : reciprocal = 16'b0000000101111010;
        8'b10101101 : reciprocal = 16'b0000000101111000;
        8'b10101110 : reciprocal = 16'b0000000101110110;
        8'b10101111 : reciprocal = 16'b0000000101110100;
        8'b10110000 : reciprocal = 16'b0000000101110010;
        8'b10110001 : reciprocal = 16'b0000000101110000;
        8'b10110010 : reciprocal = 16'b0000000101101110;
        8'b10110011 : reciprocal = 16'b0000000101101100;
        8'b10110100 : reciprocal = 16'b0000000101101010;
        8'b10110101 : reciprocal = 16'b0000000101101000;
        8'b10110110 : reciprocal = 16'b0000000101100110;
        8'b10110111 : reciprocal = 16'b0000000101100100;
        8'b10111000 : reciprocal = 16'b0000000101100010;
        8'b10111001 : reciprocal = 16'b0000000101100000;
        8'b10111010 : reciprocal = 16'b0000000101011110;
        8'b10111011 : reciprocal = 16'b0000000101011100;
        8'b10111100 : reciprocal = 16'b0000000101011010;
        8'b10111101 : reciprocal = 16'b0000000101011000;
        8'b10111110 : reciprocal = 16'b0000000101010111;
        8'b10111111 : reciprocal = 16'b0000000101010101;
        8'b11000000 : reciprocal = 16'b0000000101010011;
        8'b11000001 : reciprocal = 16'b0000000101010001;
        8'b11000010 : reciprocal = 16'b0000000101010000;
        8'b11000011 : reciprocal = 16'b0000000101001110;
        8'b11000100 : reciprocal = 16'b0000000101001100;
        8'b11000101 : reciprocal = 16'b0000000101001010;
        8'b11000110 : reciprocal = 16'b0000000101001001;
        8'b11000111 : reciprocal = 16'b0000000101000111;
        8'b11001000 : reciprocal = 16'b0000000101000110;
        8'b11001001 : reciprocal = 16'b0000000101000100;
        8'b11001010 : reciprocal = 16'b0000000101000010;
        8'b11001011 : reciprocal = 16'b0000000101000001;
        8'b11001100 : reciprocal = 16'b0000000100111111;
        8'b11001101 : reciprocal = 16'b0000000100111110;
        8'b11001110 : reciprocal = 16'b0000000100111100;
        8'b11001111 : reciprocal = 16'b0000000100111011;
        8'b11010000 : reciprocal = 16'b0000000100111001;
        8'b11010001 : reciprocal = 16'b0000000100111000;
        8'b11010010 : reciprocal = 16'b0000000100110110;
        8'b11010011 : reciprocal = 16'b0000000100110101;
        8'b11010100 : reciprocal = 16'b0000000100110011;
        8'b11010101 : reciprocal = 16'b0000000100110010;
        8'b11010110 : reciprocal = 16'b0000000100110000;
        8'b11010111 : reciprocal = 16'b0000000100101111;
        8'b11011000 : reciprocal = 16'b0000000100101110;
        8'b11011001 : reciprocal = 16'b0000000100101100;
        8'b11011010 : reciprocal = 16'b0000000100101011;
        8'b11011011 : reciprocal = 16'b0000000100101001;
        8'b11011100 : reciprocal = 16'b0000000100101000;
        8'b11011101 : reciprocal = 16'b0000000100100111;
        8'b11011110 : reciprocal = 16'b0000000100100101;
        8'b11011111 : reciprocal = 16'b0000000100100100;
        8'b11100000 : reciprocal = 16'b0000000100100011;
        8'b11100001 : reciprocal = 16'b0000000100100001;
        8'b11100010 : reciprocal = 16'b0000000100100000;
        8'b11100011 : reciprocal = 16'b0000000100011111;
        8'b11100100 : reciprocal = 16'b0000000100011110;
        8'b11100101 : reciprocal = 16'b0000000100011100;
        8'b11100110 : reciprocal = 16'b0000000100011011;
        8'b11100111 : reciprocal = 16'b0000000100011010;
        8'b11101000 : reciprocal = 16'b0000000100011001;
        8'b11101001 : reciprocal = 16'b0000000100011000;
        8'b11101010 : reciprocal = 16'b0000000100010110;
        8'b11101011 : reciprocal = 16'b0000000100010101;
        8'b11101100 : reciprocal = 16'b0000000100010100;
        8'b11101101 : reciprocal = 16'b0000000100010011;
        8'b11101110 : reciprocal = 16'b0000000100010010;
        8'b11101111 : reciprocal = 16'b0000000100010001;
        8'b11110000 : reciprocal = 16'b0000000100001111;
        8'b11110001 : reciprocal = 16'b0000000100001110;
        8'b11110010 : reciprocal = 16'b0000000100001101;
        8'b11110011 : reciprocal = 16'b0000000100001100;
        8'b11110100 : reciprocal = 16'b0000000100001011;
        8'b11110101 : reciprocal = 16'b0000000100001010;
        8'b11110110 : reciprocal = 16'b0000000100001001;
        8'b11110111 : reciprocal = 16'b0000000100001000;
        8'b11111000 : reciprocal = 16'b0000000100000111;
        8'b11111001 : reciprocal = 16'b0000000100000110;
        8'b11111010 : reciprocal = 16'b0000000100000101;
        8'b11111011 : reciprocal = 16'b0000000100000100;
        8'b11111100 : reciprocal = 16'b0000000100000011;
        8'b11111101 : reciprocal = 16'b0000000100000010;
        8'b11111110 : reciprocal = 16'b0000000100000001;
        8'b11111111 : reciprocal = 16'b0000000100000000;


        endcase
    end
    



    //////////////////////// For testbenching ////////////////////////
    // synthesis translate_off

    // synthesis translate_on

endmodule
