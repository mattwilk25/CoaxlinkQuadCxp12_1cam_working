module udivision_LUT_10bit_int_to_10bit_frac #(
)(
    input logic [10-1:0] number_in,
    output logic [10-1:0] reciprocal

);

    logic [2**10-1:0] reciprocal_LUT [10-1:0];

    always_comb begin
        case (number_in)
        10'b0000000000 : reciprocal = 10'b1111111111;
        10'b0000000001 : reciprocal = 10'b1000000000;
        10'b0000000010 : reciprocal = 10'b0101010101;
        10'b0000000011 : reciprocal = 10'b0100000000;
        10'b0000000100 : reciprocal = 10'b0011001100;
        10'b0000000101 : reciprocal = 10'b0010101010;
        10'b0000000110 : reciprocal = 10'b0010010010;
        10'b0000000111 : reciprocal = 10'b0010000000;
        10'b0000001000 : reciprocal = 10'b0001110001;
        10'b0000001001 : reciprocal = 10'b0001100110;
        10'b0000001010 : reciprocal = 10'b0001011101;
        10'b0000001011 : reciprocal = 10'b0001010101;
        10'b0000001100 : reciprocal = 10'b0001001110;
        10'b0000001101 : reciprocal = 10'b0001001001;
        10'b0000001110 : reciprocal = 10'b0001000100;
        10'b0000001111 : reciprocal = 10'b0001000000;
        10'b0000010000 : reciprocal = 10'b0000111100;
        10'b0000010001 : reciprocal = 10'b0000111000;
        10'b0000010010 : reciprocal = 10'b0000110101;
        10'b0000010011 : reciprocal = 10'b0000110011;
        10'b0000010100 : reciprocal = 10'b0000110000;
        10'b0000010101 : reciprocal = 10'b0000101110;
        10'b0000010110 : reciprocal = 10'b0000101100;
        10'b0000010111 : reciprocal = 10'b0000101010;
        10'b0000011000 : reciprocal = 10'b0000101000;
        10'b0000011001 : reciprocal = 10'b0000100111;
        10'b0000011010 : reciprocal = 10'b0000100101;
        10'b0000011011 : reciprocal = 10'b0000100100;
        10'b0000011100 : reciprocal = 10'b0000100011;
        10'b0000011101 : reciprocal = 10'b0000100010;
        10'b0000011110 : reciprocal = 10'b0000100001;
        10'b0000011111 : reciprocal = 10'b0000100000;
        10'b0000100000 : reciprocal = 10'b0000011111;
        10'b0000100001 : reciprocal = 10'b0000011110;
        10'b0000100010 : reciprocal = 10'b0000011101;
        10'b0000100011 : reciprocal = 10'b0000011100;
        10'b0000100100 : reciprocal = 10'b0000011011;
        10'b0000100101 : reciprocal = 10'b0000011010;
        10'b0000100110 : reciprocal = 10'b0000011010;
        10'b0000100111 : reciprocal = 10'b0000011001;
        10'b0000101000 : reciprocal = 10'b0000011000;
        10'b0000101001 : reciprocal = 10'b0000011000;
        10'b0000101010 : reciprocal = 10'b0000010111;
        10'b0000101011 : reciprocal = 10'b0000010111;
        10'b0000101100 : reciprocal = 10'b0000010110;
        10'b0000101101 : reciprocal = 10'b0000010110;
        10'b0000101110 : reciprocal = 10'b0000010101;
        10'b0000101111 : reciprocal = 10'b0000010101;
        10'b0000110000 : reciprocal = 10'b0000010100;
        10'b0000110001 : reciprocal = 10'b0000010100;
        10'b0000110010 : reciprocal = 10'b0000010100;
        10'b0000110011 : reciprocal = 10'b0000010011;
        10'b0000110100 : reciprocal = 10'b0000010011;
        10'b0000110101 : reciprocal = 10'b0000010010;
        10'b0000110110 : reciprocal = 10'b0000010010;
        10'b0000110111 : reciprocal = 10'b0000010010;
        10'b0000111000 : reciprocal = 10'b0000010001;
        10'b0000111001 : reciprocal = 10'b0000010001;
        10'b0000111010 : reciprocal = 10'b0000010001;
        10'b0000111011 : reciprocal = 10'b0000010001;
        10'b0000111100 : reciprocal = 10'b0000010000;
        10'b0000111101 : reciprocal = 10'b0000010000;
        10'b0000111110 : reciprocal = 10'b0000010000;
        10'b0000111111 : reciprocal = 10'b0000010000;
        10'b0001000000 : reciprocal = 10'b0000001111;
        10'b0001000001 : reciprocal = 10'b0000001111;
        10'b0001000010 : reciprocal = 10'b0000001111;
        10'b0001000011 : reciprocal = 10'b0000001111;
        10'b0001000100 : reciprocal = 10'b0000001110;
        10'b0001000101 : reciprocal = 10'b0000001110;
        10'b0001000110 : reciprocal = 10'b0000001110;
        10'b0001000111 : reciprocal = 10'b0000001110;
        10'b0001001000 : reciprocal = 10'b0000001110;
        10'b0001001001 : reciprocal = 10'b0000001101;
        10'b0001001010 : reciprocal = 10'b0000001101;
        10'b0001001011 : reciprocal = 10'b0000001101;
        10'b0001001100 : reciprocal = 10'b0000001101;
        10'b0001001101 : reciprocal = 10'b0000001101;
        10'b0001001110 : reciprocal = 10'b0000001100;
        10'b0001001111 : reciprocal = 10'b0000001100;
        10'b0001010000 : reciprocal = 10'b0000001100;
        10'b0001010001 : reciprocal = 10'b0000001100;
        10'b0001010010 : reciprocal = 10'b0000001100;
        10'b0001010011 : reciprocal = 10'b0000001100;
        10'b0001010100 : reciprocal = 10'b0000001100;
        10'b0001010101 : reciprocal = 10'b0000001011;
        10'b0001010110 : reciprocal = 10'b0000001011;
        10'b0001010111 : reciprocal = 10'b0000001011;
        10'b0001011000 : reciprocal = 10'b0000001011;
        10'b0001011001 : reciprocal = 10'b0000001011;
        10'b0001011010 : reciprocal = 10'b0000001011;
        10'b0001011011 : reciprocal = 10'b0000001011;
        10'b0001011100 : reciprocal = 10'b0000001011;
        10'b0001011101 : reciprocal = 10'b0000001010;
        10'b0001011110 : reciprocal = 10'b0000001010;
        10'b0001011111 : reciprocal = 10'b0000001010;
        10'b0001100000 : reciprocal = 10'b0000001010;
        10'b0001100001 : reciprocal = 10'b0000001010;
        10'b0001100010 : reciprocal = 10'b0000001010;
        10'b0001100011 : reciprocal = 10'b0000001010;
        10'b0001100100 : reciprocal = 10'b0000001010;
        10'b0001100101 : reciprocal = 10'b0000001010;
        10'b0001100110 : reciprocal = 10'b0000001001;
        10'b0001100111 : reciprocal = 10'b0000001001;
        10'b0001101000 : reciprocal = 10'b0000001001;
        10'b0001101001 : reciprocal = 10'b0000001001;
        10'b0001101010 : reciprocal = 10'b0000001001;
        10'b0001101011 : reciprocal = 10'b0000001001;
        10'b0001101100 : reciprocal = 10'b0000001001;
        10'b0001101101 : reciprocal = 10'b0000001001;
        10'b0001101110 : reciprocal = 10'b0000001001;
        10'b0001101111 : reciprocal = 10'b0000001001;
        10'b0001110000 : reciprocal = 10'b0000001001;
        10'b0001110001 : reciprocal = 10'b0000001000;
        10'b0001110010 : reciprocal = 10'b0000001000;
        10'b0001110011 : reciprocal = 10'b0000001000;
        10'b0001110100 : reciprocal = 10'b0000001000;
        10'b0001110101 : reciprocal = 10'b0000001000;
        10'b0001110110 : reciprocal = 10'b0000001000;
        10'b0001110111 : reciprocal = 10'b0000001000;
        10'b0001111000 : reciprocal = 10'b0000001000;
        10'b0001111001 : reciprocal = 10'b0000001000;
        10'b0001111010 : reciprocal = 10'b0000001000;
        10'b0001111011 : reciprocal = 10'b0000001000;
        10'b0001111100 : reciprocal = 10'b0000001000;
        10'b0001111101 : reciprocal = 10'b0000001000;
        10'b0001111110 : reciprocal = 10'b0000001000;
        10'b0001111111 : reciprocal = 10'b0000001000;
        10'b0010000000 : reciprocal = 10'b0000000111;
        10'b0010000001 : reciprocal = 10'b0000000111;
        10'b0010000010 : reciprocal = 10'b0000000111;
        10'b0010000011 : reciprocal = 10'b0000000111;
        10'b0010000100 : reciprocal = 10'b0000000111;
        10'b0010000101 : reciprocal = 10'b0000000111;
        10'b0010000110 : reciprocal = 10'b0000000111;
        10'b0010000111 : reciprocal = 10'b0000000111;
        10'b0010001000 : reciprocal = 10'b0000000111;
        10'b0010001001 : reciprocal = 10'b0000000111;
        10'b0010001010 : reciprocal = 10'b0000000111;
        10'b0010001011 : reciprocal = 10'b0000000111;
        10'b0010001100 : reciprocal = 10'b0000000111;
        10'b0010001101 : reciprocal = 10'b0000000111;
        10'b0010001110 : reciprocal = 10'b0000000111;
        10'b0010001111 : reciprocal = 10'b0000000111;
        10'b0010010000 : reciprocal = 10'b0000000111;
        10'b0010010001 : reciprocal = 10'b0000000111;
        10'b0010010010 : reciprocal = 10'b0000000110;
        10'b0010010011 : reciprocal = 10'b0000000110;
        10'b0010010100 : reciprocal = 10'b0000000110;
        10'b0010010101 : reciprocal = 10'b0000000110;
        10'b0010010110 : reciprocal = 10'b0000000110;
        10'b0010010111 : reciprocal = 10'b0000000110;
        10'b0010011000 : reciprocal = 10'b0000000110;
        10'b0010011001 : reciprocal = 10'b0000000110;
        10'b0010011010 : reciprocal = 10'b0000000110;
        10'b0010011011 : reciprocal = 10'b0000000110;
        10'b0010011100 : reciprocal = 10'b0000000110;
        10'b0010011101 : reciprocal = 10'b0000000110;
        10'b0010011110 : reciprocal = 10'b0000000110;
        10'b0010011111 : reciprocal = 10'b0000000110;
        10'b0010100000 : reciprocal = 10'b0000000110;
        10'b0010100001 : reciprocal = 10'b0000000110;
        10'b0010100010 : reciprocal = 10'b0000000110;
        10'b0010100011 : reciprocal = 10'b0000000110;
        10'b0010100100 : reciprocal = 10'b0000000110;
        10'b0010100101 : reciprocal = 10'b0000000110;
        10'b0010100110 : reciprocal = 10'b0000000110;
        10'b0010100111 : reciprocal = 10'b0000000110;
        10'b0010101000 : reciprocal = 10'b0000000110;
        10'b0010101001 : reciprocal = 10'b0000000110;
        10'b0010101010 : reciprocal = 10'b0000000101;
        10'b0010101011 : reciprocal = 10'b0000000101;
        10'b0010101100 : reciprocal = 10'b0000000101;
        10'b0010101101 : reciprocal = 10'b0000000101;
        10'b0010101110 : reciprocal = 10'b0000000101;
        10'b0010101111 : reciprocal = 10'b0000000101;
        10'b0010110000 : reciprocal = 10'b0000000101;
        10'b0010110001 : reciprocal = 10'b0000000101;
        10'b0010110010 : reciprocal = 10'b0000000101;
        10'b0010110011 : reciprocal = 10'b0000000101;
        10'b0010110100 : reciprocal = 10'b0000000101;
        10'b0010110101 : reciprocal = 10'b0000000101;
        10'b0010110110 : reciprocal = 10'b0000000101;
        10'b0010110111 : reciprocal = 10'b0000000101;
        10'b0010111000 : reciprocal = 10'b0000000101;
        10'b0010111001 : reciprocal = 10'b0000000101;
        10'b0010111010 : reciprocal = 10'b0000000101;
        10'b0010111011 : reciprocal = 10'b0000000101;
        10'b0010111100 : reciprocal = 10'b0000000101;
        10'b0010111101 : reciprocal = 10'b0000000101;
        10'b0010111110 : reciprocal = 10'b0000000101;
        10'b0010111111 : reciprocal = 10'b0000000101;
        10'b0011000000 : reciprocal = 10'b0000000101;
        10'b0011000001 : reciprocal = 10'b0000000101;
        10'b0011000010 : reciprocal = 10'b0000000101;
        10'b0011000011 : reciprocal = 10'b0000000101;
        10'b0011000100 : reciprocal = 10'b0000000101;
        10'b0011000101 : reciprocal = 10'b0000000101;
        10'b0011000110 : reciprocal = 10'b0000000101;
        10'b0011000111 : reciprocal = 10'b0000000101;
        10'b0011001000 : reciprocal = 10'b0000000101;
        10'b0011001001 : reciprocal = 10'b0000000101;
        10'b0011001010 : reciprocal = 10'b0000000101;
        10'b0011001011 : reciprocal = 10'b0000000101;
        10'b0011001100 : reciprocal = 10'b0000000100;
        10'b0011001101 : reciprocal = 10'b0000000100;
        10'b0011001110 : reciprocal = 10'b0000000100;
        10'b0011001111 : reciprocal = 10'b0000000100;
        10'b0011010000 : reciprocal = 10'b0000000100;
        10'b0011010001 : reciprocal = 10'b0000000100;
        10'b0011010010 : reciprocal = 10'b0000000100;
        10'b0011010011 : reciprocal = 10'b0000000100;
        10'b0011010100 : reciprocal = 10'b0000000100;
        10'b0011010101 : reciprocal = 10'b0000000100;
        10'b0011010110 : reciprocal = 10'b0000000100;
        10'b0011010111 : reciprocal = 10'b0000000100;
        10'b0011011000 : reciprocal = 10'b0000000100;
        10'b0011011001 : reciprocal = 10'b0000000100;
        10'b0011011010 : reciprocal = 10'b0000000100;
        10'b0011011011 : reciprocal = 10'b0000000100;
        10'b0011011100 : reciprocal = 10'b0000000100;
        10'b0011011101 : reciprocal = 10'b0000000100;
        10'b0011011110 : reciprocal = 10'b0000000100;
        10'b0011011111 : reciprocal = 10'b0000000100;
        10'b0011100000 : reciprocal = 10'b0000000100;
        10'b0011100001 : reciprocal = 10'b0000000100;
        10'b0011100010 : reciprocal = 10'b0000000100;
        10'b0011100011 : reciprocal = 10'b0000000100;
        10'b0011100100 : reciprocal = 10'b0000000100;
        10'b0011100101 : reciprocal = 10'b0000000100;
        10'b0011100110 : reciprocal = 10'b0000000100;
        10'b0011100111 : reciprocal = 10'b0000000100;
        10'b0011101000 : reciprocal = 10'b0000000100;
        10'b0011101001 : reciprocal = 10'b0000000100;
        10'b0011101010 : reciprocal = 10'b0000000100;
        10'b0011101011 : reciprocal = 10'b0000000100;
        10'b0011101100 : reciprocal = 10'b0000000100;
        10'b0011101101 : reciprocal = 10'b0000000100;
        10'b0011101110 : reciprocal = 10'b0000000100;
        10'b0011101111 : reciprocal = 10'b0000000100;
        10'b0011110000 : reciprocal = 10'b0000000100;
        10'b0011110001 : reciprocal = 10'b0000000100;
        10'b0011110010 : reciprocal = 10'b0000000100;
        10'b0011110011 : reciprocal = 10'b0000000100;
        10'b0011110100 : reciprocal = 10'b0000000100;
        10'b0011110101 : reciprocal = 10'b0000000100;
        10'b0011110110 : reciprocal = 10'b0000000100;
        10'b0011110111 : reciprocal = 10'b0000000100;
        10'b0011111000 : reciprocal = 10'b0000000100;
        10'b0011111001 : reciprocal = 10'b0000000100;
        10'b0011111010 : reciprocal = 10'b0000000100;
        10'b0011111011 : reciprocal = 10'b0000000100;
        10'b0011111100 : reciprocal = 10'b0000000100;
        10'b0011111101 : reciprocal = 10'b0000000100;
        10'b0011111110 : reciprocal = 10'b0000000100;
        10'b0011111111 : reciprocal = 10'b0000000100;
        10'b0100000000 : reciprocal = 10'b0000000011;
        10'b0100000001 : reciprocal = 10'b0000000011;
        10'b0100000010 : reciprocal = 10'b0000000011;
        10'b0100000011 : reciprocal = 10'b0000000011;
        10'b0100000100 : reciprocal = 10'b0000000011;
        10'b0100000101 : reciprocal = 10'b0000000011;
        10'b0100000110 : reciprocal = 10'b0000000011;
        10'b0100000111 : reciprocal = 10'b0000000011;
        10'b0100001000 : reciprocal = 10'b0000000011;
        10'b0100001001 : reciprocal = 10'b0000000011;
        10'b0100001010 : reciprocal = 10'b0000000011;
        10'b0100001011 : reciprocal = 10'b0000000011;
        10'b0100001100 : reciprocal = 10'b0000000011;
        10'b0100001101 : reciprocal = 10'b0000000011;
        10'b0100001110 : reciprocal = 10'b0000000011;
        10'b0100001111 : reciprocal = 10'b0000000011;
        10'b0100010000 : reciprocal = 10'b0000000011;
        10'b0100010001 : reciprocal = 10'b0000000011;
        10'b0100010010 : reciprocal = 10'b0000000011;
        10'b0100010011 : reciprocal = 10'b0000000011;
        10'b0100010100 : reciprocal = 10'b0000000011;
        10'b0100010101 : reciprocal = 10'b0000000011;
        10'b0100010110 : reciprocal = 10'b0000000011;
        10'b0100010111 : reciprocal = 10'b0000000011;
        10'b0100011000 : reciprocal = 10'b0000000011;
        10'b0100011001 : reciprocal = 10'b0000000011;
        10'b0100011010 : reciprocal = 10'b0000000011;
        10'b0100011011 : reciprocal = 10'b0000000011;
        10'b0100011100 : reciprocal = 10'b0000000011;
        10'b0100011101 : reciprocal = 10'b0000000011;
        10'b0100011110 : reciprocal = 10'b0000000011;
        10'b0100011111 : reciprocal = 10'b0000000011;
        10'b0100100000 : reciprocal = 10'b0000000011;
        10'b0100100001 : reciprocal = 10'b0000000011;
        10'b0100100010 : reciprocal = 10'b0000000011;
        10'b0100100011 : reciprocal = 10'b0000000011;
        10'b0100100100 : reciprocal = 10'b0000000011;
        10'b0100100101 : reciprocal = 10'b0000000011;
        10'b0100100110 : reciprocal = 10'b0000000011;
        10'b0100100111 : reciprocal = 10'b0000000011;
        10'b0100101000 : reciprocal = 10'b0000000011;
        10'b0100101001 : reciprocal = 10'b0000000011;
        10'b0100101010 : reciprocal = 10'b0000000011;
        10'b0100101011 : reciprocal = 10'b0000000011;
        10'b0100101100 : reciprocal = 10'b0000000011;
        10'b0100101101 : reciprocal = 10'b0000000011;
        10'b0100101110 : reciprocal = 10'b0000000011;
        10'b0100101111 : reciprocal = 10'b0000000011;
        10'b0100110000 : reciprocal = 10'b0000000011;
        10'b0100110001 : reciprocal = 10'b0000000011;
        10'b0100110010 : reciprocal = 10'b0000000011;
        10'b0100110011 : reciprocal = 10'b0000000011;
        10'b0100110100 : reciprocal = 10'b0000000011;
        10'b0100110101 : reciprocal = 10'b0000000011;
        10'b0100110110 : reciprocal = 10'b0000000011;
        10'b0100110111 : reciprocal = 10'b0000000011;
        10'b0100111000 : reciprocal = 10'b0000000011;
        10'b0100111001 : reciprocal = 10'b0000000011;
        10'b0100111010 : reciprocal = 10'b0000000011;
        10'b0100111011 : reciprocal = 10'b0000000011;
        10'b0100111100 : reciprocal = 10'b0000000011;
        10'b0100111101 : reciprocal = 10'b0000000011;
        10'b0100111110 : reciprocal = 10'b0000000011;
        10'b0100111111 : reciprocal = 10'b0000000011;
        10'b0101000000 : reciprocal = 10'b0000000011;
        10'b0101000001 : reciprocal = 10'b0000000011;
        10'b0101000010 : reciprocal = 10'b0000000011;
        10'b0101000011 : reciprocal = 10'b0000000011;
        10'b0101000100 : reciprocal = 10'b0000000011;
        10'b0101000101 : reciprocal = 10'b0000000011;
        10'b0101000110 : reciprocal = 10'b0000000011;
        10'b0101000111 : reciprocal = 10'b0000000011;
        10'b0101001000 : reciprocal = 10'b0000000011;
        10'b0101001001 : reciprocal = 10'b0000000011;
        10'b0101001010 : reciprocal = 10'b0000000011;
        10'b0101001011 : reciprocal = 10'b0000000011;
        10'b0101001100 : reciprocal = 10'b0000000011;
        10'b0101001101 : reciprocal = 10'b0000000011;
        10'b0101001110 : reciprocal = 10'b0000000011;
        10'b0101001111 : reciprocal = 10'b0000000011;
        10'b0101010000 : reciprocal = 10'b0000000011;
        10'b0101010001 : reciprocal = 10'b0000000011;
        10'b0101010010 : reciprocal = 10'b0000000011;
        10'b0101010011 : reciprocal = 10'b0000000011;
        10'b0101010100 : reciprocal = 10'b0000000011;
        10'b0101010101 : reciprocal = 10'b0000000010;
        10'b0101010110 : reciprocal = 10'b0000000010;
        10'b0101010111 : reciprocal = 10'b0000000010;
        10'b0101011000 : reciprocal = 10'b0000000010;
        10'b0101011001 : reciprocal = 10'b0000000010;
        10'b0101011010 : reciprocal = 10'b0000000010;
        10'b0101011011 : reciprocal = 10'b0000000010;
        10'b0101011100 : reciprocal = 10'b0000000010;
        10'b0101011101 : reciprocal = 10'b0000000010;
        10'b0101011110 : reciprocal = 10'b0000000010;
        10'b0101011111 : reciprocal = 10'b0000000010;
        10'b0101100000 : reciprocal = 10'b0000000010;
        10'b0101100001 : reciprocal = 10'b0000000010;
        10'b0101100010 : reciprocal = 10'b0000000010;
        10'b0101100011 : reciprocal = 10'b0000000010;
        10'b0101100100 : reciprocal = 10'b0000000010;
        10'b0101100101 : reciprocal = 10'b0000000010;
        10'b0101100110 : reciprocal = 10'b0000000010;
        10'b0101100111 : reciprocal = 10'b0000000010;
        10'b0101101000 : reciprocal = 10'b0000000010;
        10'b0101101001 : reciprocal = 10'b0000000010;
        10'b0101101010 : reciprocal = 10'b0000000010;
        10'b0101101011 : reciprocal = 10'b0000000010;
        10'b0101101100 : reciprocal = 10'b0000000010;
        10'b0101101101 : reciprocal = 10'b0000000010;
        10'b0101101110 : reciprocal = 10'b0000000010;
        10'b0101101111 : reciprocal = 10'b0000000010;
        10'b0101110000 : reciprocal = 10'b0000000010;
        10'b0101110001 : reciprocal = 10'b0000000010;
        10'b0101110010 : reciprocal = 10'b0000000010;
        10'b0101110011 : reciprocal = 10'b0000000010;
        10'b0101110100 : reciprocal = 10'b0000000010;
        10'b0101110101 : reciprocal = 10'b0000000010;
        10'b0101110110 : reciprocal = 10'b0000000010;
        10'b0101110111 : reciprocal = 10'b0000000010;
        10'b0101111000 : reciprocal = 10'b0000000010;
        10'b0101111001 : reciprocal = 10'b0000000010;
        10'b0101111010 : reciprocal = 10'b0000000010;
        10'b0101111011 : reciprocal = 10'b0000000010;
        10'b0101111100 : reciprocal = 10'b0000000010;
        10'b0101111101 : reciprocal = 10'b0000000010;
        10'b0101111110 : reciprocal = 10'b0000000010;
        10'b0101111111 : reciprocal = 10'b0000000010;
        10'b0110000000 : reciprocal = 10'b0000000010;
        10'b0110000001 : reciprocal = 10'b0000000010;
        10'b0110000010 : reciprocal = 10'b0000000010;
        10'b0110000011 : reciprocal = 10'b0000000010;
        10'b0110000100 : reciprocal = 10'b0000000010;
        10'b0110000101 : reciprocal = 10'b0000000010;
        10'b0110000110 : reciprocal = 10'b0000000010;
        10'b0110000111 : reciprocal = 10'b0000000010;
        10'b0110001000 : reciprocal = 10'b0000000010;
        10'b0110001001 : reciprocal = 10'b0000000010;
        10'b0110001010 : reciprocal = 10'b0000000010;
        10'b0110001011 : reciprocal = 10'b0000000010;
        10'b0110001100 : reciprocal = 10'b0000000010;
        10'b0110001101 : reciprocal = 10'b0000000010;
        10'b0110001110 : reciprocal = 10'b0000000010;
        10'b0110001111 : reciprocal = 10'b0000000010;
        10'b0110010000 : reciprocal = 10'b0000000010;
        10'b0110010001 : reciprocal = 10'b0000000010;
        10'b0110010010 : reciprocal = 10'b0000000010;
        10'b0110010011 : reciprocal = 10'b0000000010;
        10'b0110010100 : reciprocal = 10'b0000000010;
        10'b0110010101 : reciprocal = 10'b0000000010;
        10'b0110010110 : reciprocal = 10'b0000000010;
        10'b0110010111 : reciprocal = 10'b0000000010;
        10'b0110011000 : reciprocal = 10'b0000000010;
        10'b0110011001 : reciprocal = 10'b0000000010;
        10'b0110011010 : reciprocal = 10'b0000000010;
        10'b0110011011 : reciprocal = 10'b0000000010;
        10'b0110011100 : reciprocal = 10'b0000000010;
        10'b0110011101 : reciprocal = 10'b0000000010;
        10'b0110011110 : reciprocal = 10'b0000000010;
        10'b0110011111 : reciprocal = 10'b0000000010;
        10'b0110100000 : reciprocal = 10'b0000000010;
        10'b0110100001 : reciprocal = 10'b0000000010;
        10'b0110100010 : reciprocal = 10'b0000000010;
        10'b0110100011 : reciprocal = 10'b0000000010;
        10'b0110100100 : reciprocal = 10'b0000000010;
        10'b0110100101 : reciprocal = 10'b0000000010;
        10'b0110100110 : reciprocal = 10'b0000000010;
        10'b0110100111 : reciprocal = 10'b0000000010;
        10'b0110101000 : reciprocal = 10'b0000000010;
        10'b0110101001 : reciprocal = 10'b0000000010;
        10'b0110101010 : reciprocal = 10'b0000000010;
        10'b0110101011 : reciprocal = 10'b0000000010;
        10'b0110101100 : reciprocal = 10'b0000000010;
        10'b0110101101 : reciprocal = 10'b0000000010;
        10'b0110101110 : reciprocal = 10'b0000000010;
        10'b0110101111 : reciprocal = 10'b0000000010;
        10'b0110110000 : reciprocal = 10'b0000000010;
        10'b0110110001 : reciprocal = 10'b0000000010;
        10'b0110110010 : reciprocal = 10'b0000000010;
        10'b0110110011 : reciprocal = 10'b0000000010;
        10'b0110110100 : reciprocal = 10'b0000000010;
        10'b0110110101 : reciprocal = 10'b0000000010;
        10'b0110110110 : reciprocal = 10'b0000000010;
        10'b0110110111 : reciprocal = 10'b0000000010;
        10'b0110111000 : reciprocal = 10'b0000000010;
        10'b0110111001 : reciprocal = 10'b0000000010;
        10'b0110111010 : reciprocal = 10'b0000000010;
        10'b0110111011 : reciprocal = 10'b0000000010;
        10'b0110111100 : reciprocal = 10'b0000000010;
        10'b0110111101 : reciprocal = 10'b0000000010;
        10'b0110111110 : reciprocal = 10'b0000000010;
        10'b0110111111 : reciprocal = 10'b0000000010;
        10'b0111000000 : reciprocal = 10'b0000000010;
        10'b0111000001 : reciprocal = 10'b0000000010;
        10'b0111000010 : reciprocal = 10'b0000000010;
        10'b0111000011 : reciprocal = 10'b0000000010;
        10'b0111000100 : reciprocal = 10'b0000000010;
        10'b0111000101 : reciprocal = 10'b0000000010;
        10'b0111000110 : reciprocal = 10'b0000000010;
        10'b0111000111 : reciprocal = 10'b0000000010;
        10'b0111001000 : reciprocal = 10'b0000000010;
        10'b0111001001 : reciprocal = 10'b0000000010;
        10'b0111001010 : reciprocal = 10'b0000000010;
        10'b0111001011 : reciprocal = 10'b0000000010;
        10'b0111001100 : reciprocal = 10'b0000000010;
        10'b0111001101 : reciprocal = 10'b0000000010;
        10'b0111001110 : reciprocal = 10'b0000000010;
        10'b0111001111 : reciprocal = 10'b0000000010;
        10'b0111010000 : reciprocal = 10'b0000000010;
        10'b0111010001 : reciprocal = 10'b0000000010;
        10'b0111010010 : reciprocal = 10'b0000000010;
        10'b0111010011 : reciprocal = 10'b0000000010;
        10'b0111010100 : reciprocal = 10'b0000000010;
        10'b0111010101 : reciprocal = 10'b0000000010;
        10'b0111010110 : reciprocal = 10'b0000000010;
        10'b0111010111 : reciprocal = 10'b0000000010;
        10'b0111011000 : reciprocal = 10'b0000000010;
        10'b0111011001 : reciprocal = 10'b0000000010;
        10'b0111011010 : reciprocal = 10'b0000000010;
        10'b0111011011 : reciprocal = 10'b0000000010;
        10'b0111011100 : reciprocal = 10'b0000000010;
        10'b0111011101 : reciprocal = 10'b0000000010;
        10'b0111011110 : reciprocal = 10'b0000000010;
        10'b0111011111 : reciprocal = 10'b0000000010;
        10'b0111100000 : reciprocal = 10'b0000000010;
        10'b0111100001 : reciprocal = 10'b0000000010;
        10'b0111100010 : reciprocal = 10'b0000000010;
        10'b0111100011 : reciprocal = 10'b0000000010;
        10'b0111100100 : reciprocal = 10'b0000000010;
        10'b0111100101 : reciprocal = 10'b0000000010;
        10'b0111100110 : reciprocal = 10'b0000000010;
        10'b0111100111 : reciprocal = 10'b0000000010;
        10'b0111101000 : reciprocal = 10'b0000000010;
        10'b0111101001 : reciprocal = 10'b0000000010;
        10'b0111101010 : reciprocal = 10'b0000000010;
        10'b0111101011 : reciprocal = 10'b0000000010;
        10'b0111101100 : reciprocal = 10'b0000000010;
        10'b0111101101 : reciprocal = 10'b0000000010;
        10'b0111101110 : reciprocal = 10'b0000000010;
        10'b0111101111 : reciprocal = 10'b0000000010;
        10'b0111110000 : reciprocal = 10'b0000000010;
        10'b0111110001 : reciprocal = 10'b0000000010;
        10'b0111110010 : reciprocal = 10'b0000000010;
        10'b0111110011 : reciprocal = 10'b0000000010;
        10'b0111110100 : reciprocal = 10'b0000000010;
        10'b0111110101 : reciprocal = 10'b0000000010;
        10'b0111110110 : reciprocal = 10'b0000000010;
        10'b0111110111 : reciprocal = 10'b0000000010;
        10'b0111111000 : reciprocal = 10'b0000000010;
        10'b0111111001 : reciprocal = 10'b0000000010;
        10'b0111111010 : reciprocal = 10'b0000000010;
        10'b0111111011 : reciprocal = 10'b0000000010;
        10'b0111111100 : reciprocal = 10'b0000000010;
        10'b0111111101 : reciprocal = 10'b0000000010;
        10'b0111111110 : reciprocal = 10'b0000000010;
        10'b0111111111 : reciprocal = 10'b0000000010;
        default : reciprocal = 10'b0000000001;


        endcase
    end
    



    //////////////////////// For testbenching ////////////////////////
    // synthesis translate_off

    // synthesis translate_on

endmodule
