module udivision_LUT_8bit_int_to_32bit_frac #(
)(
    input logic [8-1:0] number_in,
    output logic [32-1:0] reciprocal

);

    logic [2**8-1:0] reciprocal_LUT [32-1:0];

    always_comb begin
        case (number_in)
        8'b00000000 : reciprocal = 32'b11111111111111111111111111111111;
        8'b00000001 : reciprocal = 32'b10000000000000000000000000000000;
        8'b00000010 : reciprocal = 32'b01010101010101010101010101010101;
        8'b00000011 : reciprocal = 32'b01000000000000000000000000000000;
        8'b00000100 : reciprocal = 32'b00110011001100110011001100110011;
        8'b00000101 : reciprocal = 32'b00101010101010101010101010101010;
        8'b00000110 : reciprocal = 32'b00100100100100100100100100100100;
        8'b00000111 : reciprocal = 32'b00100000000000000000000000000000;
        8'b00001000 : reciprocal = 32'b00011100011100011100011100011100;
        8'b00001001 : reciprocal = 32'b00011001100110011001100110011001;
        8'b00001010 : reciprocal = 32'b00010111010001011101000101110100;
        8'b00001011 : reciprocal = 32'b00010101010101010101010101010101;
        8'b00001100 : reciprocal = 32'b00010011101100010011101100010011;
        8'b00001101 : reciprocal = 32'b00010010010010010010010010010010;
        8'b00001110 : reciprocal = 32'b00010001000100010001000100010001;
        8'b00001111 : reciprocal = 32'b00010000000000000000000000000000;
        8'b00010000 : reciprocal = 32'b00001111000011110000111100001111;
        8'b00010001 : reciprocal = 32'b00001110001110001110001110001110;
        8'b00010010 : reciprocal = 32'b00001101011110010100001101011110;
        8'b00010011 : reciprocal = 32'b00001100110011001100110011001100;
        8'b00010100 : reciprocal = 32'b00001100001100001100001100001100;
        8'b00010101 : reciprocal = 32'b00001011101000101110100010111010;
        8'b00010110 : reciprocal = 32'b00001011001000010110010000101100;
        8'b00010111 : reciprocal = 32'b00001010101010101010101010101010;
        8'b00011000 : reciprocal = 32'b00001010001111010111000010100011;
        8'b00011001 : reciprocal = 32'b00001001110110001001110110001001;
        8'b00011010 : reciprocal = 32'b00001001011110110100001001011110;
        8'b00011011 : reciprocal = 32'b00001001001001001001001001001001;
        8'b00011100 : reciprocal = 32'b00001000110100111101110010110000;
        8'b00011101 : reciprocal = 32'b00001000100010001000100010001000;
        8'b00011110 : reciprocal = 32'b00001000010000100001000010000100;
        8'b00011111 : reciprocal = 32'b00001000000000000000000000000000;
        8'b00100000 : reciprocal = 32'b00000111110000011111000001111100;
        8'b00100001 : reciprocal = 32'b00000111100001111000011110000111;
        8'b00100010 : reciprocal = 32'b00000111010100000111010100000111;
        8'b00100011 : reciprocal = 32'b00000111000111000111000111000111;
        8'b00100100 : reciprocal = 32'b00000110111010110011111001000101;
        8'b00100101 : reciprocal = 32'b00000110101111001010000110101111;
        8'b00100110 : reciprocal = 32'b00000110100100000110100100000110;
        8'b00100111 : reciprocal = 32'b00000110011001100110011001100110;
        8'b00101000 : reciprocal = 32'b00000110001111100111000001100011;
        8'b00101001 : reciprocal = 32'b00000110000110000110000110000110;
        8'b00101010 : reciprocal = 32'b00000101111101000001011111010000;
        8'b00101011 : reciprocal = 32'b00000101110100010111010001011101;
        8'b00101100 : reciprocal = 32'b00000101101100000101101100000101;
        8'b00101101 : reciprocal = 32'b00000101100100001011001000010110;
        8'b00101110 : reciprocal = 32'b00000101011100100110001000001010;
        8'b00101111 : reciprocal = 32'b00000101010101010101010101010101;
        8'b00110000 : reciprocal = 32'b00000101001110010111100000101001;
        8'b00110001 : reciprocal = 32'b00000101000111101011100001010001;
        8'b00110010 : reciprocal = 32'b00000101000001010000010100000101;
        8'b00110011 : reciprocal = 32'b00000100111011000100111011000100;
        8'b00110100 : reciprocal = 32'b00000100110101001000011100111110;
        8'b00110101 : reciprocal = 32'b00000100101111011010000100101111;
        8'b00110110 : reciprocal = 32'b00000100101001111001000001001010;
        8'b00110111 : reciprocal = 32'b00000100100100100100100100100100;
        8'b00111000 : reciprocal = 32'b00000100011111011100000100011111;
        8'b00111001 : reciprocal = 32'b00000100011010011110111001011000;
        8'b00111010 : reciprocal = 32'b00000100010101101100011110010111;
        8'b00111011 : reciprocal = 32'b00000100010001000100010001000100;
        8'b00111100 : reciprocal = 32'b00000100001100100101110001010011;
        8'b00111101 : reciprocal = 32'b00000100001000010000100001000010;
        8'b00111110 : reciprocal = 32'b00000100000100000100000100000100;
        8'b00111111 : reciprocal = 32'b00000100000000000000000000000000;
        8'b01000000 : reciprocal = 32'b00000011111100000011111100000011;
        8'b01000001 : reciprocal = 32'b00000011111000001111100000111110;
        8'b01000010 : reciprocal = 32'b00000011110100100010011000110101;
        8'b01000011 : reciprocal = 32'b00000011110000111100001111000011;
        8'b01000100 : reciprocal = 32'b00000011101101011100110000001110;
        8'b01000101 : reciprocal = 32'b00000011101010000011101010000011;
        8'b01000110 : reciprocal = 32'b00000011100110110000101011010001;
        8'b01000111 : reciprocal = 32'b00000011100011100011100011100011;
        8'b01001000 : reciprocal = 32'b00000011100000011100000011100000;
        8'b01001001 : reciprocal = 32'b00000011011101011001111100100010;
        8'b01001010 : reciprocal = 32'b00000011011010011101000000110110;
        8'b01001011 : reciprocal = 32'b00000011010111100101000011010111;
        8'b01001100 : reciprocal = 32'b00000011010100110001110111101100;
        8'b01001101 : reciprocal = 32'b00000011010010000011010010000011;
        8'b01001110 : reciprocal = 32'b00000011001111011001000111010010;
        8'b01001111 : reciprocal = 32'b00000011001100110011001100110011;
        8'b01010000 : reciprocal = 32'b00000011001010010001011000011111;
        8'b01010001 : reciprocal = 32'b00000011000111110011100000110001;
        8'b01010010 : reciprocal = 32'b00000011000101011001011100100001;
        8'b01010011 : reciprocal = 32'b00000011000011000011000011000011;
        8'b01010100 : reciprocal = 32'b00000011000000110000001100000011;
        8'b01010101 : reciprocal = 32'b00000010111110100000101111101000;
        8'b01010110 : reciprocal = 32'b00000010111100010100100110010000;
        8'b01010111 : reciprocal = 32'b00000010111010001011101000101110;
        8'b01011000 : reciprocal = 32'b00000010111000000101110000001011;
        8'b01011001 : reciprocal = 32'b00000010110110000010110110000010;
        8'b01011010 : reciprocal = 32'b00000010110100000010110100000010;
        8'b01011011 : reciprocal = 32'b00000010110010000101100100001011;
        8'b01011100 : reciprocal = 32'b00000010110000001011000000101100;
        8'b01011101 : reciprocal = 32'b00000010101110010011000100000101;
        8'b01011110 : reciprocal = 32'b00000010101100011101101001000110;
        8'b01011111 : reciprocal = 32'b00000010101010101010101010101010;
        8'b01100000 : reciprocal = 32'b00000010101000111010000011111101;
        8'b01100001 : reciprocal = 32'b00000010100111001011110000010100;
        8'b01100010 : reciprocal = 32'b00000010100101011111101011010100;
        8'b01100011 : reciprocal = 32'b00000010100011110101110000101000;
        8'b01100100 : reciprocal = 32'b00000010100010001101111100001100;
        8'b01100101 : reciprocal = 32'b00000010100000101000001010000010;
        8'b01100110 : reciprocal = 32'b00000010011111000100010110010111;
        8'b01100111 : reciprocal = 32'b00000010011101100010011101100010;
        8'b01101000 : reciprocal = 32'b00000010011100000010011100000010;
        8'b01101001 : reciprocal = 32'b00000010011010100100001110011111;
        8'b01101010 : reciprocal = 32'b00000010011001000111110001101001;
        8'b01101011 : reciprocal = 32'b00000010010111101101000010010111;
        8'b01101100 : reciprocal = 32'b00000010010110010011111101101001;
        8'b01101101 : reciprocal = 32'b00000010010100111100100000100101;
        8'b01101110 : reciprocal = 32'b00000010010011100110101000010111;
        8'b01101111 : reciprocal = 32'b00000010010010010010010010010010;
        8'b01110000 : reciprocal = 32'b00000010010000111111011011110000;
        8'b01110001 : reciprocal = 32'b00000010001111101110000010001111;
        8'b01110010 : reciprocal = 32'b00000010001110011110000011010101;
        8'b01110011 : reciprocal = 32'b00000010001101001111011100101100;
        8'b01110100 : reciprocal = 32'b00000010001100000010001100000010;
        8'b01110101 : reciprocal = 32'b00000010001010110110001111001011;
        8'b01110110 : reciprocal = 32'b00000010001001101011100100000010;
        8'b01110111 : reciprocal = 32'b00000010001000100010001000100010;
        8'b01111000 : reciprocal = 32'b00000010000111011001111010101101;
        8'b01111001 : reciprocal = 32'b00000010000110010010111000101001;
        8'b01111010 : reciprocal = 32'b00000010000101001101000000100001;
        8'b01111011 : reciprocal = 32'b00000010000100001000010000100001;
        8'b01111100 : reciprocal = 32'b00000010000011000100100110111010;
        8'b01111101 : reciprocal = 32'b00000010000010000010000010000010;
        8'b01111110 : reciprocal = 32'b00000010000001000000100000010000;
        8'b01111111 : reciprocal = 32'b00000010000000000000000000000000;
        8'b10000000 : reciprocal = 32'b00000001111111000000011111110000;
        8'b10000001 : reciprocal = 32'b00000001111110000001111110000001;
        8'b10000010 : reciprocal = 32'b00000001111101000100011001011001;
        8'b10000011 : reciprocal = 32'b00000001111100000111110000011111;
        8'b10000100 : reciprocal = 32'b00000001111011001100000001111011;
        8'b10000101 : reciprocal = 32'b00000001111010010001001100011010;
        8'b10000110 : reciprocal = 32'b00000001111001010111001110101100;
        8'b10000111 : reciprocal = 32'b00000001111000011110000111100001;
        8'b10001000 : reciprocal = 32'b00000001110111100101110101101110;
        8'b10001001 : reciprocal = 32'b00000001110110101110011000000111;
        8'b10001010 : reciprocal = 32'b00000001110101110111101101100101;
        8'b10001011 : reciprocal = 32'b00000001110101000001110101000001;
        8'b10001100 : reciprocal = 32'b00000001110100001100101101011000;
        8'b10001101 : reciprocal = 32'b00000001110011011000010101101000;
        8'b10001110 : reciprocal = 32'b00000001110010100100101100110000;
        8'b10001111 : reciprocal = 32'b00000001110001110001110001110001;
        8'b10010000 : reciprocal = 32'b00000001110000111111100011110000;
        8'b10010001 : reciprocal = 32'b00000001110000001110000001110000;
        8'b10010010 : reciprocal = 32'b00000001101111011101001010111000;
        8'b10010011 : reciprocal = 32'b00000001101110101100111110010001;
        8'b10010100 : reciprocal = 32'b00000001101101111101011011000011;
        8'b10010101 : reciprocal = 32'b00000001101101001110100000011011;
        8'b10010110 : reciprocal = 32'b00000001101100100000001101100100;
        8'b10010111 : reciprocal = 32'b00000001101011110010100001101011;
        8'b10011000 : reciprocal = 32'b00000001101011000101011100000001;
        8'b10011001 : reciprocal = 32'b00000001101010011000111011110110;
        8'b10011010 : reciprocal = 32'b00000001101001101101000000011010;
        8'b10011011 : reciprocal = 32'b00000001101001000001101001000001;
        8'b10011100 : reciprocal = 32'b00000001101000010110110100111111;
        8'b10011101 : reciprocal = 32'b00000001100111101100100011101001;
        8'b10011110 : reciprocal = 32'b00000001100111000010110100010100;
        8'b10011111 : reciprocal = 32'b00000001100110011001100110011001;
        8'b10100000 : reciprocal = 32'b00000001100101110000111001001111;
        8'b10100001 : reciprocal = 32'b00000001100101001000101100001111;
        8'b10100010 : reciprocal = 32'b00000001100100100000111110110100;
        8'b10100011 : reciprocal = 32'b00000001100011111001110000011000;
        8'b10100100 : reciprocal = 32'b00000001100011010011000000011000;
        8'b10100101 : reciprocal = 32'b00000001100010101100101110010000;
        8'b10100110 : reciprocal = 32'b00000001100010000110111001011111;
        8'b10100111 : reciprocal = 32'b00000001100001100001100001100001;
        8'b10101000 : reciprocal = 32'b00000001100000111100100101110111;
        8'b10101001 : reciprocal = 32'b00000001100000011000000110000001;
        8'b10101010 : reciprocal = 32'b00000001011111110100000001011111;
        8'b10101011 : reciprocal = 32'b00000001011111010000010111110100;
        8'b10101100 : reciprocal = 32'b00000001011110101101001000100000;
        8'b10101101 : reciprocal = 32'b00000001011110001010010011001000;
        8'b10101110 : reciprocal = 32'b00000001011101100111110111001110;
        8'b10101111 : reciprocal = 32'b00000001011101000101110100010111;
        8'b10110000 : reciprocal = 32'b00000001011100100100001010000111;
        8'b10110001 : reciprocal = 32'b00000001011100000010111000000101;
        8'b10110010 : reciprocal = 32'b00000001011011100001111101110110;
        8'b10110011 : reciprocal = 32'b00000001011011000001011011000001;
        8'b10110100 : reciprocal = 32'b00000001011010100001001111001101;
        8'b10110101 : reciprocal = 32'b00000001011010000001011010000001;
        8'b10110110 : reciprocal = 32'b00000001011001100001111011000110;
        8'b10110111 : reciprocal = 32'b00000001011001000010110010000101;
        8'b10111000 : reciprocal = 32'b00000001011000100011111110100111;
        8'b10111001 : reciprocal = 32'b00000001011000000101100000010110;
        8'b10111010 : reciprocal = 32'b00000001010111100111010110111011;
        8'b10111011 : reciprocal = 32'b00000001010111001001100010000010;
        8'b10111100 : reciprocal = 32'b00000001010110101100000001010110;
        8'b10111101 : reciprocal = 32'b00000001010110001110110100100011;
        8'b10111110 : reciprocal = 32'b00000001010101110001111011010011;
        8'b10111111 : reciprocal = 32'b00000001010101010101010101010101;
        8'b11000000 : reciprocal = 32'b00000001010100111001000010010100;
        8'b11000001 : reciprocal = 32'b00000001010100011101000001111110;
        8'b11000010 : reciprocal = 32'b00000001010100000001010100000001;
        8'b11000011 : reciprocal = 32'b00000001010011100101111000001010;
        8'b11000100 : reciprocal = 32'b00000001010011001010101110001000;
        8'b11000101 : reciprocal = 32'b00000001010010101111110101101010;
        8'b11000110 : reciprocal = 32'b00000001010010010101001110011110;
        8'b11000111 : reciprocal = 32'b00000001010001111010111000010100;
        8'b11001000 : reciprocal = 32'b00000001010001100000110010111100;
        8'b11001001 : reciprocal = 32'b00000001010001000110111110000110;
        8'b11001010 : reciprocal = 32'b00000001010000101101011001100010;
        8'b11001011 : reciprocal = 32'b00000001010000010100000101000001;
        8'b11001100 : reciprocal = 32'b00000001001111111011000000010011;
        8'b11001101 : reciprocal = 32'b00000001001111100010001011001011;
        8'b11001110 : reciprocal = 32'b00000001001111001001100101011010;
        8'b11001111 : reciprocal = 32'b00000001001110110001001110110001;
        8'b11010000 : reciprocal = 32'b00000001001110011001000111000010;
        8'b11010001 : reciprocal = 32'b00000001001110000001001110000001;
        8'b11010010 : reciprocal = 32'b00000001001101101001100011011111;
        8'b11010011 : reciprocal = 32'b00000001001101010010000111001111;
        8'b11010100 : reciprocal = 32'b00000001001100111010111001000101;
        8'b11010101 : reciprocal = 32'b00000001001100100011111000110100;
        8'b11010110 : reciprocal = 32'b00000001001100001101000110010000;
        8'b11010111 : reciprocal = 32'b00000001001011110110100001001011;
        8'b11011000 : reciprocal = 32'b00000001001011100000001001011100;
        8'b11011001 : reciprocal = 32'b00000001001011001001111110110100;
        8'b11011010 : reciprocal = 32'b00000001001010110100000001001010;
        8'b11011011 : reciprocal = 32'b00000001001010011110010000010010;
        8'b11011100 : reciprocal = 32'b00000001001010001000101100000001;
        8'b11011101 : reciprocal = 32'b00000001001001110011010100001011;
        8'b11011110 : reciprocal = 32'b00000001001001011110001000100111;
        8'b11011111 : reciprocal = 32'b00000001001001001001001001001001;
        8'b11100000 : reciprocal = 32'b00000001001000110100010101100111;
        8'b11100001 : reciprocal = 32'b00000001001000011111101101111000;
        8'b11100010 : reciprocal = 32'b00000001001000001011010001110000;
        8'b11100011 : reciprocal = 32'b00000001000111110111000001000111;
        8'b11100100 : reciprocal = 32'b00000001000111100010111011110011;
        8'b11100101 : reciprocal = 32'b00000001000111001111000001101010;
        8'b11100110 : reciprocal = 32'b00000001000110111011010010100100;
        8'b11100111 : reciprocal = 32'b00000001000110100111101110010110;
        8'b11101000 : reciprocal = 32'b00000001000110010100010100111000;
        8'b11101001 : reciprocal = 32'b00000001000110000001000110000001;
        8'b11101010 : reciprocal = 32'b00000001000101101110000001101000;
        8'b11101011 : reciprocal = 32'b00000001000101011011000111100101;
        8'b11101100 : reciprocal = 32'b00000001000101001000010111110000;
        8'b11101101 : reciprocal = 32'b00000001000100110101110010000001;
        8'b11101110 : reciprocal = 32'b00000001000100100011010110001110;
        8'b11101111 : reciprocal = 32'b00000001000100010001000100010001;
        8'b11110000 : reciprocal = 32'b00000001000011111110111100000001;
        8'b11110001 : reciprocal = 32'b00000001000011101100111101010110;
        8'b11110010 : reciprocal = 32'b00000001000011011011001000001010;
        8'b11110011 : reciprocal = 32'b00000001000011001001011100010100;
        8'b11110100 : reciprocal = 32'b00000001000010110111111001101110;
        8'b11110101 : reciprocal = 32'b00000001000010100110100000010000;
        8'b11110110 : reciprocal = 32'b00000001000010010101001111110011;
        8'b11110111 : reciprocal = 32'b00000001000010000100001000010000;
        8'b11111000 : reciprocal = 32'b00000001000001110011001001100000;
        8'b11111001 : reciprocal = 32'b00000001000001100010010011011101;
        8'b11111010 : reciprocal = 32'b00000001000001010001100101111111;
        8'b11111011 : reciprocal = 32'b00000001000001000001000001000001;
        8'b11111100 : reciprocal = 32'b00000001000000110000100100011011;
        8'b11111101 : reciprocal = 32'b00000001000000100000010000001000;
        8'b11111110 : reciprocal = 32'b00000001000000010000000100000001;
        8'b11111111 : reciprocal = 32'b00000001000000000000000000000000;


        endcase
    end
    



    //////////////////////// For testbenching ////////////////////////
    // synthesis translate_off

    // synthesis translate_on

endmodule
